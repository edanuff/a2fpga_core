// Generated build timestamp
`define BUILD_DATETIME "20250808154519"
