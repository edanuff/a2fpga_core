// Generated build timestamp
`define BUILD_DATETIME "20250808010411"
