`define CONSOLE_60K
