// Generated build timestamp
`define BUILD_DATETIME "20250827083518"
